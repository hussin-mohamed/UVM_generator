module sva (
    //variables
);
//assertions 
    endmodule